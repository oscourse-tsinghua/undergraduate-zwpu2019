// pico_cyc10_qys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module pico_cyc10_qys (
		input  wire       clk_clk,       //   clk.clk
		output wire [7:0] led_export,    //   led.export
		input  wire       reset_reset_n, // reset.reset_n
		output wire [7:0] seg_export,    //   seg.export
		output wire       trap_export,   //  trap.export
		input  wire       uart_rxd,      //  uart.rxd
		output wire       uart_txd       //      .txd
	);

	wire  [31:0] pico_cyc10_0_altera_axi4lite_master_awaddr;  // pico_cyc10_0:axm_awaddr -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_awaddr
	wire   [1:0] pico_cyc10_0_altera_axi4lite_master_bresp;   // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_bresp -> pico_cyc10_0:axm_bresp
	wire         pico_cyc10_0_altera_axi4lite_master_arready; // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_arready -> pico_cyc10_0:axm_arready
	wire  [31:0] pico_cyc10_0_altera_axi4lite_master_rdata;   // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_rdata -> pico_cyc10_0:axm_rdata
	wire         pico_cyc10_0_altera_axi4lite_master_wready;  // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_wready -> pico_cyc10_0:axm_wready
	wire   [3:0] pico_cyc10_0_altera_axi4lite_master_wstrb;   // pico_cyc10_0:axm_wstrb -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_wstrb
	wire         pico_cyc10_0_altera_axi4lite_master_awready; // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_awready -> pico_cyc10_0:axm_awready
	wire         pico_cyc10_0_altera_axi4lite_master_rready;  // pico_cyc10_0:axm_rready -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_rready
	wire         pico_cyc10_0_altera_axi4lite_master_bready;  // pico_cyc10_0:axm_bready -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_bready
	wire         pico_cyc10_0_altera_axi4lite_master_wvalid;  // pico_cyc10_0:axm_wvalid -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_wvalid
	wire  [31:0] pico_cyc10_0_altera_axi4lite_master_araddr;  // pico_cyc10_0:axm_araddr -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_araddr
	wire   [2:0] pico_cyc10_0_altera_axi4lite_master_arprot;  // pico_cyc10_0:axm_arprot -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_arprot
	wire   [1:0] pico_cyc10_0_altera_axi4lite_master_rresp;   // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_rresp -> pico_cyc10_0:axm_rresp
	wire   [2:0] pico_cyc10_0_altera_axi4lite_master_awprot;  // pico_cyc10_0:axm_awprot -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_awprot
	wire  [31:0] pico_cyc10_0_altera_axi4lite_master_wdata;   // pico_cyc10_0:axm_wdata -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_wdata
	wire         pico_cyc10_0_altera_axi4lite_master_arvalid; // pico_cyc10_0:axm_arvalid -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_arvalid
	wire         pico_cyc10_0_altera_axi4lite_master_bvalid;  // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_bvalid -> pico_cyc10_0:axm_bvalid
	wire         pico_cyc10_0_altera_axi4lite_master_awvalid; // pico_cyc10_0:axm_awvalid -> mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_awvalid
	wire         pico_cyc10_0_altera_axi4lite_master_rvalid;  // mm_interconnect_0:pico_cyc10_0_altera_axi4lite_master_rvalid -> pico_cyc10_0:axm_rvalid
	wire         mm_interconnect_0_rom_s1_chipselect;         // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;           // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;        // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire  [13:0] mm_interconnect_0_rom_s1_address;            // mm_interconnect_0:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;         // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_0_rom_s1_write;              // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;          // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_0_rom_s1_clken;              // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         mm_interconnect_0_ram_s1_chipselect;         // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;           // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;            // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;         // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;              // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;          // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;              // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_led_s1_chipselect;         // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;           // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;            // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;              // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;          // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_seg_s1_chipselect;         // mm_interconnect_0:seg_s1_chipselect -> seg:chipselect
	wire  [31:0] mm_interconnect_0_seg_s1_readdata;           // seg:readdata -> mm_interconnect_0:seg_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_s1_address;            // mm_interconnect_0:seg_s1_address -> seg:address
	wire         mm_interconnect_0_seg_s1_write;              // mm_interconnect_0:seg_s1_write -> seg:write_n
	wire  [31:0] mm_interconnect_0_seg_s1_writedata;          // mm_interconnect_0:seg_s1_writedata -> seg:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;      // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;        // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;         // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;            // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;   // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;           // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;       // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         irq_mapper_receiver0_irq;                    // uart_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] pico_cyc10_0_interrupt_receiver_0_irq;       // irq_mapper:sender_irq -> pico_cyc10_0:inr_irq
	wire         rst_controller_reset_out_reset;              // rst_controller:reset_out -> [irq_mapper:reset, led:reset_n, mm_interconnect_0:pico_cyc10_0_reset_reset_bridge_in_reset_reset, pico_cyc10_0:rsi_resetn, ram:reset, rom:reset, rst_translator:in_reset, seg:reset_n, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;          // rst_controller:reset_req -> [ram:reset_req, rom:reset_req, rst_translator:reset_req_in]

	pico_cyc10_qys_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	picorv32_axi_wrapper #(
		.ENABLE_COUNTERS      (2'b01),
		.ENABLE_COUNTERS64    (2'b01),
		.ENABLE_REGS_16_31    (2'b01),
		.ENABLE_REGS_DUALPORT (2'b01),
		.TWO_STAGE_SHIFT      (2'b01),
		.BARREL_SHIFTER       (2'b00),
		.TWO_CYCLE_COMPARE    (2'b00),
		.TWO_CYCLE_ALU        (2'b00),
		.COMPRESSED_ISA       (2'b00),
		.CATCH_MISALIGN       (2'b01),
		.CATCH_ILLINSN        (2'b01),
		.ENABLE_PCPI          (2'b00),
		.ENABLE_MUL           (2'b01),
		.ENABLE_FAST_MUL      (2'b00),
		.ENABLE_DIV           (2'b01),
		.ENABLE_IRQ           (2'b01),
		.ENABLE_IRQ_QREGS     (2'b01),
		.ENABLE_IRQ_TIMER     (2'b01),
		.ENABLE_TRACE         (2'b00),
		.REGS_INIT_ZERO       (2'b00),
		.MASKED_IRQ           (34'b0000000000000000000000000000000000),
		.LATCHED_IRQ          (34'b0011111111111111111111111111111111),
		.PROGADDR_RESET       (34'b0000000000000000000000000000000000),
		.PROGADDR_IRQ         (34'b0000000000000000000000000000010000),
		.STACKADDR            (34'b0011111111111111111111111111111111)
	) pico_cyc10_0 (
		.clk         (clk_clk),                                     //                  clock.clk
		.rsi_resetn  (~rst_controller_reset_out_reset),             //                  reset.reset_n
		.coe_trap    (trap_export),                                 //          conduit_end_0.export
		.inr_irq     (pico_cyc10_0_interrupt_receiver_0_irq),       //   interrupt_receiver_0.irq
		.axm_awvalid (pico_cyc10_0_altera_axi4lite_master_awvalid), // altera_axi4lite_master.awvalid
		.axm_awready (pico_cyc10_0_altera_axi4lite_master_awready), //                       .awready
		.axm_awaddr  (pico_cyc10_0_altera_axi4lite_master_awaddr),  //                       .awaddr
		.axm_awprot  (pico_cyc10_0_altera_axi4lite_master_awprot),  //                       .awprot
		.axm_wvalid  (pico_cyc10_0_altera_axi4lite_master_wvalid),  //                       .wvalid
		.axm_wready  (pico_cyc10_0_altera_axi4lite_master_wready),  //                       .wready
		.axm_wdata   (pico_cyc10_0_altera_axi4lite_master_wdata),   //                       .wdata
		.axm_wstrb   (pico_cyc10_0_altera_axi4lite_master_wstrb),   //                       .wstrb
		.axm_bvalid  (pico_cyc10_0_altera_axi4lite_master_bvalid),  //                       .bvalid
		.axm_bresp   (pico_cyc10_0_altera_axi4lite_master_bresp),   //                       .bresp
		.axm_bready  (pico_cyc10_0_altera_axi4lite_master_bready),  //                       .bready
		.axm_arvalid (pico_cyc10_0_altera_axi4lite_master_arvalid), //                       .arvalid
		.axm_arready (pico_cyc10_0_altera_axi4lite_master_arready), //                       .arready
		.axm_araddr  (pico_cyc10_0_altera_axi4lite_master_araddr),  //                       .araddr
		.axm_arprot  (pico_cyc10_0_altera_axi4lite_master_arprot),  //                       .arprot
		.axm_rvalid  (pico_cyc10_0_altera_axi4lite_master_rvalid),  //                       .rvalid
		.axm_rresp   (pico_cyc10_0_altera_axi4lite_master_rresp),   //                       .rresp
		.axm_rready  (pico_cyc10_0_altera_axi4lite_master_rready),  //                       .rready
		.axm_rdata   (pico_cyc10_0_altera_axi4lite_master_rdata)    //                       .rdata
	);

	pico_cyc10_qys_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	pico_cyc10_qys_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	pico_cyc10_qys_seg seg (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_s1_readdata),   //                    .readdata
		.out_port   (seg_export)                           // external_connection.export
	);

	pico_cyc10_qys_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                  // external_connection.export
		.txd           (uart_txd),                                  //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	pico_cyc10_qys_mm_interconnect_0 mm_interconnect_0 (
		.pico_cyc10_0_altera_axi4lite_master_awaddr     (pico_cyc10_0_altera_axi4lite_master_awaddr),  //      pico_cyc10_0_altera_axi4lite_master.awaddr
		.pico_cyc10_0_altera_axi4lite_master_awprot     (pico_cyc10_0_altera_axi4lite_master_awprot),  //                                         .awprot
		.pico_cyc10_0_altera_axi4lite_master_awvalid    (pico_cyc10_0_altera_axi4lite_master_awvalid), //                                         .awvalid
		.pico_cyc10_0_altera_axi4lite_master_awready    (pico_cyc10_0_altera_axi4lite_master_awready), //                                         .awready
		.pico_cyc10_0_altera_axi4lite_master_wdata      (pico_cyc10_0_altera_axi4lite_master_wdata),   //                                         .wdata
		.pico_cyc10_0_altera_axi4lite_master_wstrb      (pico_cyc10_0_altera_axi4lite_master_wstrb),   //                                         .wstrb
		.pico_cyc10_0_altera_axi4lite_master_wvalid     (pico_cyc10_0_altera_axi4lite_master_wvalid),  //                                         .wvalid
		.pico_cyc10_0_altera_axi4lite_master_wready     (pico_cyc10_0_altera_axi4lite_master_wready),  //                                         .wready
		.pico_cyc10_0_altera_axi4lite_master_bresp      (pico_cyc10_0_altera_axi4lite_master_bresp),   //                                         .bresp
		.pico_cyc10_0_altera_axi4lite_master_bvalid     (pico_cyc10_0_altera_axi4lite_master_bvalid),  //                                         .bvalid
		.pico_cyc10_0_altera_axi4lite_master_bready     (pico_cyc10_0_altera_axi4lite_master_bready),  //                                         .bready
		.pico_cyc10_0_altera_axi4lite_master_araddr     (pico_cyc10_0_altera_axi4lite_master_araddr),  //                                         .araddr
		.pico_cyc10_0_altera_axi4lite_master_arprot     (pico_cyc10_0_altera_axi4lite_master_arprot),  //                                         .arprot
		.pico_cyc10_0_altera_axi4lite_master_arvalid    (pico_cyc10_0_altera_axi4lite_master_arvalid), //                                         .arvalid
		.pico_cyc10_0_altera_axi4lite_master_arready    (pico_cyc10_0_altera_axi4lite_master_arready), //                                         .arready
		.pico_cyc10_0_altera_axi4lite_master_rdata      (pico_cyc10_0_altera_axi4lite_master_rdata),   //                                         .rdata
		.pico_cyc10_0_altera_axi4lite_master_rresp      (pico_cyc10_0_altera_axi4lite_master_rresp),   //                                         .rresp
		.pico_cyc10_0_altera_axi4lite_master_rvalid     (pico_cyc10_0_altera_axi4lite_master_rvalid),  //                                         .rvalid
		.pico_cyc10_0_altera_axi4lite_master_rready     (pico_cyc10_0_altera_axi4lite_master_rready),  //                                         .rready
		.clk_0_clk_clk                                  (clk_clk),                                     //                                clk_0_clk.clk
		.pico_cyc10_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),              // pico_cyc10_0_reset_reset_bridge_in_reset.reset
		.led_s1_address                                 (mm_interconnect_0_led_s1_address),            //                                   led_s1.address
		.led_s1_write                                   (mm_interconnect_0_led_s1_write),              //                                         .write
		.led_s1_readdata                                (mm_interconnect_0_led_s1_readdata),           //                                         .readdata
		.led_s1_writedata                               (mm_interconnect_0_led_s1_writedata),          //                                         .writedata
		.led_s1_chipselect                              (mm_interconnect_0_led_s1_chipselect),         //                                         .chipselect
		.ram_s1_address                                 (mm_interconnect_0_ram_s1_address),            //                                   ram_s1.address
		.ram_s1_write                                   (mm_interconnect_0_ram_s1_write),              //                                         .write
		.ram_s1_readdata                                (mm_interconnect_0_ram_s1_readdata),           //                                         .readdata
		.ram_s1_writedata                               (mm_interconnect_0_ram_s1_writedata),          //                                         .writedata
		.ram_s1_byteenable                              (mm_interconnect_0_ram_s1_byteenable),         //                                         .byteenable
		.ram_s1_chipselect                              (mm_interconnect_0_ram_s1_chipselect),         //                                         .chipselect
		.ram_s1_clken                                   (mm_interconnect_0_ram_s1_clken),              //                                         .clken
		.rom_s1_address                                 (mm_interconnect_0_rom_s1_address),            //                                   rom_s1.address
		.rom_s1_write                                   (mm_interconnect_0_rom_s1_write),              //                                         .write
		.rom_s1_readdata                                (mm_interconnect_0_rom_s1_readdata),           //                                         .readdata
		.rom_s1_writedata                               (mm_interconnect_0_rom_s1_writedata),          //                                         .writedata
		.rom_s1_byteenable                              (mm_interconnect_0_rom_s1_byteenable),         //                                         .byteenable
		.rom_s1_chipselect                              (mm_interconnect_0_rom_s1_chipselect),         //                                         .chipselect
		.rom_s1_clken                                   (mm_interconnect_0_rom_s1_clken),              //                                         .clken
		.rom_s1_debugaccess                             (mm_interconnect_0_rom_s1_debugaccess),        //                                         .debugaccess
		.seg_s1_address                                 (mm_interconnect_0_seg_s1_address),            //                                   seg_s1.address
		.seg_s1_write                                   (mm_interconnect_0_seg_s1_write),              //                                         .write
		.seg_s1_readdata                                (mm_interconnect_0_seg_s1_readdata),           //                                         .readdata
		.seg_s1_writedata                               (mm_interconnect_0_seg_s1_writedata),          //                                         .writedata
		.seg_s1_chipselect                              (mm_interconnect_0_seg_s1_chipselect),         //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),         //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),           //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),            //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),        //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),       //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),   //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)       //                                         .chipselect
	);

	pico_cyc10_qys_irq_mapper irq_mapper (
		.clk           (clk_clk),                               //       clk.clk
		.reset         (rst_controller_reset_out_reset),        // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),              // receiver0.irq
		.sender_irq    (pico_cyc10_0_interrupt_receiver_0_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
